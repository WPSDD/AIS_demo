library verilog;
use verilog.vl_types.all;
entity tb_dehdlc is
end tb_dehdlc;
