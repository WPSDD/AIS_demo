library verilog;
use verilog.vl_types.all;
entity tb_pad_test is
end tb_pad_test;
