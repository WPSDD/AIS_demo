library verilog;
use verilog.vl_types.all;
entity tb_dds_18M is
end tb_dds_18M;
