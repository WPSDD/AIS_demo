library verilog;
use verilog.vl_types.all;
entity tb_denrzi is
end tb_denrzi;
